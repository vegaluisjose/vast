module one_param # (
    parameter width = 32)(
    input wire [3:0] data);
endmodule