module bar ();
endmodule