module module_with_always_comb ();
    always_comb begin
        $display("hello world");
    end
endmodule
