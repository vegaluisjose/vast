module two_params # (
    parameter width = 4,
    parameter length = 8)(
    input wire [3:0] data);
endmodule