module foo ();
endmodule