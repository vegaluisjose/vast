module one_input (
    input wire [4:0] a);
endmodule