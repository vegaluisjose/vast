module module_with_initial ();
    initial begin
        $display("initial");
    end
endmodule
