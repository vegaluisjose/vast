module module_with_final ();
    final begin
        $display("final");
    end
endmodule
