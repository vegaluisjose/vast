module two_params # (
    parameter width = 32'd4,
    parameter length = 32'd8)(
    input wire [3:0] data);
endmodule