module empty ();
endmodule