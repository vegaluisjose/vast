module four_inputs (
    input logic [1:0] a,
    input logic [6:0] b,
    input logic [3:0] c,
    input logic d);
endmodule