module one_wire ();
    wire [7:0] one_wire;
endmodule
