module one_input (
    input logic [4:0] a);
endmodule