module one_param # (
    parameter width = 32'd32)(
    input wire [3:0] data);
endmodule