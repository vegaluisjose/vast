module mix_params # (
    parameter width = 4,
    parameter length = 8,
    parameter name = "foo")(
    input wire [3:0] data);
endmodule