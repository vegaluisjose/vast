module three_inputs (
    input wire [4:0] a,
    input wire [60:0] b,
    input wire c);
endmodule
