module main ();
    always_comb begin
        foo(2, x);
    end
endmodule
