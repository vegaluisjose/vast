module module_with_instance_attribute ();
    (*LOC = "X0Y0", TYPE = "LUT6"*)
    prim i0 (
        .port_a(4'h0)
    );
endmodule
