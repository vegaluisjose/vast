(*use = "yes"*)
module attribute ();
endmodule
