module prim # (
    parameter WIDTH = 32'd4,
    parameter name = "foo")(
    input logic [3:0] port_a);
endmodule
